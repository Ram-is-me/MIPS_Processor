module branch_pc(in_pc,imm,branch_pc)